magic
tech sky130A
timestamp 1742229583
<< nwell >>
rect -200 -200 1600 220
rect -205 -1240 1595 -830
<< nmos >>
rect -60 -400 -45 -300
rect 190 -400 205 -300
rect 440 -400 455 -300
rect 690 -400 705 -300
rect 940 -400 955 -300
rect 1190 -400 1205 -300
rect 1440 -400 1455 -300
rect -60 -730 -45 -630
rect 190 -730 205 -630
rect 440 -730 455 -630
rect 690 -730 705 -630
rect 940 -730 955 -630
rect 1190 -730 1205 -630
rect 1440 -730 1455 -630
<< pmos >>
rect -60 -150 -45 50
rect 190 -150 205 50
rect 440 -150 455 50
rect 690 -150 705 50
rect 940 -150 955 50
rect 1190 -150 1205 50
rect 1440 -150 1455 50
rect -60 -1080 -45 -880
rect 190 -1080 205 -880
rect 440 -1080 455 -880
rect 690 -1080 705 -880
rect 940 -1080 955 -880
rect 1190 -1080 1205 -880
rect 1440 -1080 1455 -880
<< ndiff >>
rect -105 -340 -60 -300
rect -105 -360 -95 -340
rect -75 -360 -60 -340
rect -105 -400 -60 -360
rect -45 -340 0 -300
rect -45 -360 -30 -340
rect -10 -360 0 -340
rect -45 -400 0 -360
rect 145 -340 190 -300
rect 145 -360 155 -340
rect 175 -360 190 -340
rect 145 -400 190 -360
rect 205 -340 250 -300
rect 205 -360 220 -340
rect 240 -360 250 -340
rect 205 -400 250 -360
rect 395 -340 440 -300
rect 395 -360 405 -340
rect 425 -360 440 -340
rect 395 -400 440 -360
rect 455 -340 500 -300
rect 455 -360 470 -340
rect 490 -360 500 -340
rect 455 -400 500 -360
rect 645 -340 690 -300
rect 645 -360 655 -340
rect 675 -360 690 -340
rect 645 -400 690 -360
rect 705 -340 750 -300
rect 705 -360 720 -340
rect 740 -360 750 -340
rect 705 -400 750 -360
rect 895 -340 940 -300
rect 895 -360 905 -340
rect 925 -360 940 -340
rect 895 -400 940 -360
rect 955 -340 1000 -300
rect 955 -360 970 -340
rect 990 -360 1000 -340
rect 955 -400 1000 -360
rect 1145 -340 1190 -300
rect 1145 -360 1155 -340
rect 1175 -360 1190 -340
rect 1145 -400 1190 -360
rect 1205 -340 1250 -300
rect 1205 -360 1220 -340
rect 1240 -360 1250 -340
rect 1205 -400 1250 -360
rect 1395 -340 1440 -300
rect 1395 -360 1405 -340
rect 1425 -360 1440 -340
rect 1395 -400 1440 -360
rect 1455 -340 1500 -300
rect 1455 -360 1470 -340
rect 1490 -360 1500 -340
rect 1455 -400 1500 -360
rect -105 -670 -60 -630
rect -105 -690 -95 -670
rect -75 -690 -60 -670
rect -105 -730 -60 -690
rect -45 -670 0 -630
rect -45 -690 -30 -670
rect -10 -690 0 -670
rect -45 -730 0 -690
rect 145 -670 190 -630
rect 145 -690 155 -670
rect 175 -690 190 -670
rect 145 -730 190 -690
rect 205 -670 250 -630
rect 205 -690 220 -670
rect 240 -690 250 -670
rect 205 -730 250 -690
rect 395 -670 440 -630
rect 395 -690 405 -670
rect 425 -690 440 -670
rect 395 -730 440 -690
rect 455 -670 500 -630
rect 455 -690 470 -670
rect 490 -690 500 -670
rect 455 -730 500 -690
rect 645 -670 690 -630
rect 645 -690 655 -670
rect 675 -690 690 -670
rect 645 -730 690 -690
rect 705 -670 750 -630
rect 705 -690 720 -670
rect 740 -690 750 -670
rect 705 -730 750 -690
rect 895 -670 940 -630
rect 895 -690 905 -670
rect 925 -690 940 -670
rect 895 -730 940 -690
rect 955 -670 1000 -630
rect 955 -690 970 -670
rect 990 -690 1000 -670
rect 955 -730 1000 -690
rect 1145 -670 1190 -630
rect 1145 -690 1155 -670
rect 1175 -690 1190 -670
rect 1145 -730 1190 -690
rect 1205 -670 1250 -630
rect 1205 -690 1220 -670
rect 1240 -690 1250 -670
rect 1205 -730 1250 -690
rect 1395 -670 1440 -630
rect 1395 -690 1405 -670
rect 1425 -690 1440 -670
rect 1395 -730 1440 -690
rect 1455 -670 1500 -630
rect 1455 -690 1470 -670
rect 1490 -690 1500 -670
rect 1455 -730 1500 -690
<< pdiff >>
rect -105 -40 -60 50
rect -105 -60 -95 -40
rect -75 -60 -60 -40
rect -105 -150 -60 -60
rect -45 -40 0 50
rect -45 -60 -30 -40
rect -10 -60 0 -40
rect -45 -150 0 -60
rect 145 -40 190 50
rect 145 -60 155 -40
rect 175 -60 190 -40
rect 145 -150 190 -60
rect 205 -40 250 50
rect 205 -60 220 -40
rect 240 -60 250 -40
rect 205 -150 250 -60
rect 395 -40 440 50
rect 395 -60 405 -40
rect 425 -60 440 -40
rect 395 -150 440 -60
rect 455 -40 500 50
rect 455 -60 470 -40
rect 490 -60 500 -40
rect 455 -150 500 -60
rect 645 -40 690 50
rect 645 -60 655 -40
rect 675 -60 690 -40
rect 645 -150 690 -60
rect 705 -40 750 50
rect 705 -60 720 -40
rect 740 -60 750 -40
rect 705 -150 750 -60
rect 895 -40 940 50
rect 895 -60 905 -40
rect 925 -60 940 -40
rect 895 -150 940 -60
rect 955 -40 1000 50
rect 955 -60 970 -40
rect 990 -60 1000 -40
rect 955 -150 1000 -60
rect 1145 -40 1190 50
rect 1145 -60 1155 -40
rect 1175 -60 1190 -40
rect 1145 -150 1190 -60
rect 1205 -40 1250 50
rect 1205 -60 1220 -40
rect 1240 -60 1250 -40
rect 1205 -150 1250 -60
rect 1395 -40 1440 50
rect 1395 -60 1405 -40
rect 1425 -60 1440 -40
rect 1395 -150 1440 -60
rect 1455 -40 1500 50
rect 1455 -60 1470 -40
rect 1490 -60 1500 -40
rect 1455 -150 1500 -60
rect -105 -970 -60 -880
rect -105 -990 -95 -970
rect -75 -990 -60 -970
rect -105 -1080 -60 -990
rect -45 -970 0 -880
rect -45 -990 -30 -970
rect -10 -990 0 -970
rect -45 -1080 0 -990
rect 145 -970 190 -880
rect 145 -990 155 -970
rect 175 -990 190 -970
rect 145 -1080 190 -990
rect 205 -970 250 -880
rect 205 -990 220 -970
rect 240 -990 250 -970
rect 205 -1080 250 -990
rect 395 -970 440 -880
rect 395 -990 405 -970
rect 425 -990 440 -970
rect 395 -1080 440 -990
rect 455 -970 500 -880
rect 455 -990 470 -970
rect 490 -990 500 -970
rect 455 -1080 500 -990
rect 645 -970 690 -880
rect 645 -990 655 -970
rect 675 -990 690 -970
rect 645 -1080 690 -990
rect 705 -970 750 -880
rect 705 -990 720 -970
rect 740 -990 750 -970
rect 705 -1080 750 -990
rect 895 -970 940 -880
rect 895 -990 905 -970
rect 925 -990 940 -970
rect 895 -1080 940 -990
rect 955 -970 1000 -880
rect 955 -990 970 -970
rect 990 -990 1000 -970
rect 955 -1080 1000 -990
rect 1145 -970 1190 -880
rect 1145 -990 1155 -970
rect 1175 -990 1190 -970
rect 1145 -1080 1190 -990
rect 1205 -970 1250 -880
rect 1205 -990 1220 -970
rect 1240 -990 1250 -970
rect 1205 -1080 1250 -990
rect 1395 -970 1440 -880
rect 1395 -990 1405 -970
rect 1425 -990 1440 -970
rect 1395 -1080 1440 -990
rect 1455 -970 1500 -880
rect 1455 -990 1470 -970
rect 1490 -990 1500 -970
rect 1455 -1080 1500 -990
<< ndiffc >>
rect -95 -360 -75 -340
rect -30 -360 -10 -340
rect 155 -360 175 -340
rect 220 -360 240 -340
rect 405 -360 425 -340
rect 470 -360 490 -340
rect 655 -360 675 -340
rect 720 -360 740 -340
rect 905 -360 925 -340
rect 970 -360 990 -340
rect 1155 -360 1175 -340
rect 1220 -360 1240 -340
rect 1405 -360 1425 -340
rect 1470 -360 1490 -340
rect -95 -690 -75 -670
rect -30 -690 -10 -670
rect 155 -690 175 -670
rect 220 -690 240 -670
rect 405 -690 425 -670
rect 470 -690 490 -670
rect 655 -690 675 -670
rect 720 -690 740 -670
rect 905 -690 925 -670
rect 970 -690 990 -670
rect 1155 -690 1175 -670
rect 1220 -690 1240 -670
rect 1405 -690 1425 -670
rect 1470 -690 1490 -670
<< pdiffc >>
rect -95 -60 -75 -40
rect -30 -60 -10 -40
rect 155 -60 175 -40
rect 220 -60 240 -40
rect 405 -60 425 -40
rect 470 -60 490 -40
rect 655 -60 675 -40
rect 720 -60 740 -40
rect 905 -60 925 -40
rect 970 -60 990 -40
rect 1155 -60 1175 -40
rect 1220 -60 1240 -40
rect 1405 -60 1425 -40
rect 1470 -60 1490 -40
rect -95 -990 -75 -970
rect -30 -990 -10 -970
rect 155 -990 175 -970
rect 220 -990 240 -970
rect 405 -990 425 -970
rect 470 -990 490 -970
rect 655 -990 675 -970
rect 720 -990 740 -970
rect 905 -990 925 -970
rect 970 -990 990 -970
rect 1155 -990 1175 -970
rect 1220 -990 1240 -970
rect 1405 -990 1425 -970
rect 1470 -990 1490 -970
<< psubdiff >>
rect -105 -515 0 -465
rect 145 -515 250 -465
rect 395 -515 500 -465
rect 645 -515 750 -465
rect 895 -515 1000 -465
rect 1145 -515 1250 -465
rect 1395 -515 1500 -465
<< nsubdiff >>
rect -105 115 0 165
rect 145 115 250 165
rect 395 115 500 165
rect 645 115 750 165
rect 895 115 1000 165
rect 1145 115 1250 165
rect 1395 115 1500 165
rect -105 -1190 0 -1140
rect 145 -1190 250 -1140
rect 395 -1190 500 -1140
rect 645 -1190 750 -1140
rect 895 -1190 1000 -1140
rect 1145 -1190 1250 -1140
rect 1395 -1190 1500 -1140
<< poly >>
rect -60 50 -45 65
rect 190 50 205 65
rect 440 50 455 65
rect 690 50 705 65
rect 940 50 955 65
rect 1190 50 1205 65
rect 1440 50 1455 65
rect -60 -300 -45 -150
rect 190 -300 205 -150
rect 440 -300 455 -150
rect 690 -300 705 -150
rect 940 -300 955 -150
rect 1190 -170 1205 -150
rect 1440 -170 1455 -150
rect 1130 -180 1205 -170
rect 1130 -200 1140 -180
rect 1160 -200 1205 -180
rect 1130 -210 1205 -200
rect 1380 -180 1455 -170
rect 1380 -200 1390 -180
rect 1410 -200 1455 -180
rect 1380 -210 1455 -200
rect 1190 -300 1205 -210
rect 1440 -300 1455 -210
rect -60 -415 -45 -400
rect 190 -415 205 -400
rect 440 -415 455 -400
rect 690 -415 705 -400
rect 940 -415 955 -400
rect 1190 -415 1205 -400
rect 1440 -415 1455 -400
rect -60 -630 -45 -615
rect 190 -630 205 -615
rect 440 -630 455 -615
rect 690 -630 705 -615
rect 940 -630 955 -615
rect 1190 -630 1205 -615
rect 1440 -630 1455 -615
rect -60 -880 -45 -730
rect 190 -880 205 -730
rect 440 -880 455 -730
rect 690 -880 705 -730
rect 940 -880 955 -730
rect 1190 -880 1205 -730
rect 1440 -880 1455 -730
rect -60 -1095 -45 -1080
rect 190 -1095 205 -1080
rect 440 -1095 455 -1080
rect 690 -1095 705 -1080
rect 940 -1095 955 -1080
rect 1190 -1095 1205 -1080
rect 1440 -1095 1455 -1080
<< polycont >>
rect 1140 -200 1160 -180
rect 1390 -200 1410 -180
<< locali >>
rect -105 155 0 165
rect -105 125 -95 155
rect -65 125 -40 155
rect -10 125 0 155
rect -105 115 0 125
rect 145 155 250 165
rect 145 125 155 155
rect 185 125 210 155
rect 240 125 250 155
rect 145 115 250 125
rect 395 155 500 165
rect 395 125 405 155
rect 435 125 460 155
rect 490 125 500 155
rect 395 115 500 125
rect 645 155 750 165
rect 645 125 655 155
rect 685 125 710 155
rect 740 125 750 155
rect 645 115 750 125
rect 895 155 1000 165
rect 895 125 905 155
rect 935 125 960 155
rect 990 125 1000 155
rect 895 115 1000 125
rect 1145 155 1250 165
rect 1145 125 1155 155
rect 1185 125 1210 155
rect 1240 125 1250 155
rect 1145 115 1250 125
rect 1395 155 1500 165
rect 1395 125 1405 155
rect 1435 125 1460 155
rect 1490 125 1500 155
rect 1395 115 1500 125
rect -105 -40 -65 115
rect 585 70 750 90
rect -105 -60 -95 -40
rect -75 -60 -65 -40
rect -105 -150 -65 -60
rect -40 -40 0 50
rect 145 -40 185 50
rect -40 -60 -30 -40
rect -10 -60 155 -40
rect 175 -60 185 -40
rect -40 -150 0 -60
rect 145 -150 185 -60
rect 210 -40 250 50
rect 395 -40 435 50
rect 210 -60 220 -40
rect 240 -60 405 -40
rect 425 -60 435 -40
rect 210 -150 250 -60
rect 395 -150 435 -60
rect 460 -40 500 50
rect 585 -40 605 70
rect 730 50 750 70
rect 460 -60 470 -40
rect 490 -60 605 -40
rect 645 -40 685 50
rect 645 -60 655 -40
rect 675 -60 685 -40
rect 460 -150 500 -60
rect 255 -235 295 -185
rect 255 -255 265 -235
rect 285 -255 295 -235
rect 255 -260 295 -255
rect 545 -260 565 -60
rect 645 -150 685 -60
rect 710 -40 750 50
rect 710 -60 720 -40
rect 740 -60 750 -40
rect 710 -150 750 -60
rect 895 -40 935 115
rect 895 -60 905 -40
rect 925 -60 935 -40
rect 895 -150 935 -60
rect 960 -40 1000 50
rect 960 -60 970 -40
rect 990 -60 1000 -40
rect 960 -150 1000 -60
rect 1145 -40 1185 115
rect 1145 -60 1155 -40
rect 1175 -60 1185 -40
rect 1145 -150 1185 -60
rect 1210 -40 1250 50
rect 1210 -60 1220 -40
rect 1240 -60 1250 -40
rect 655 -170 675 -150
rect 970 -170 990 -150
rect 655 -190 990 -170
rect 1130 -180 1180 -170
rect 1130 -200 1140 -180
rect 1160 -200 1180 -180
rect 1130 -210 1180 -200
rect 1210 -245 1250 -60
rect 1395 -40 1435 115
rect 1395 -60 1405 -40
rect 1425 -60 1435 -40
rect 1395 -150 1435 -60
rect 1460 -40 1500 50
rect 1460 -60 1470 -40
rect 1490 -60 1500 -40
rect 1460 -165 1500 -60
rect 1380 -180 1430 -170
rect 1380 -200 1390 -180
rect 1410 -200 1430 -180
rect 1380 -210 1430 -200
rect 1460 -185 1475 -165
rect 1495 -185 1500 -165
rect 220 -280 740 -260
rect 220 -300 240 -280
rect 470 -300 490 -280
rect 720 -300 740 -280
rect 815 -280 990 -260
rect -105 -340 -65 -300
rect -105 -360 -95 -340
rect -75 -360 -65 -340
rect -105 -465 -65 -360
rect -40 -340 0 -300
rect 145 -340 185 -300
rect -40 -360 -30 -340
rect -10 -360 155 -340
rect 175 -360 185 -340
rect -40 -400 0 -360
rect 145 -400 185 -360
rect 210 -340 250 -300
rect 210 -360 220 -340
rect 240 -360 250 -340
rect 210 -400 250 -360
rect 395 -340 435 -300
rect 395 -360 405 -340
rect 425 -360 435 -340
rect 395 -400 435 -360
rect 460 -340 500 -300
rect 460 -360 470 -340
rect 490 -360 500 -340
rect 460 -400 500 -360
rect 645 -340 685 -300
rect 645 -360 655 -340
rect 675 -360 685 -340
rect 645 -400 685 -360
rect 710 -340 750 -300
rect 710 -360 720 -340
rect 740 -360 750 -340
rect 710 -400 750 -360
rect 405 -420 425 -400
rect 655 -420 675 -400
rect 815 -420 835 -280
rect 970 -300 990 -280
rect 1210 -265 1225 -245
rect 1245 -265 1250 -245
rect 405 -440 835 -420
rect 895 -340 935 -300
rect 895 -360 905 -340
rect 925 -360 935 -340
rect 895 -465 935 -360
rect 960 -340 1000 -300
rect 960 -360 970 -340
rect 990 -360 1000 -340
rect 960 -400 1000 -360
rect 1145 -340 1185 -300
rect 1145 -360 1155 -340
rect 1175 -360 1185 -340
rect 1145 -465 1185 -360
rect 1210 -340 1250 -265
rect 1210 -360 1220 -340
rect 1240 -360 1250 -340
rect 1210 -400 1250 -360
rect 1395 -340 1435 -300
rect 1395 -360 1405 -340
rect 1425 -360 1435 -340
rect 1395 -465 1435 -360
rect 1460 -340 1500 -185
rect 1460 -360 1470 -340
rect 1490 -360 1500 -340
rect 1460 -400 1500 -360
rect -105 -475 0 -465
rect -105 -505 -95 -475
rect -65 -505 -40 -475
rect -10 -505 0 -475
rect -105 -515 0 -505
rect 145 -475 250 -465
rect 145 -505 155 -475
rect 185 -505 210 -475
rect 240 -505 250 -475
rect 145 -515 250 -505
rect 395 -475 500 -465
rect 395 -505 405 -475
rect 435 -505 460 -475
rect 490 -505 500 -475
rect 395 -515 500 -505
rect 645 -475 750 -465
rect 645 -505 655 -475
rect 685 -505 710 -475
rect 740 -505 750 -475
rect 645 -515 750 -505
rect 895 -475 1000 -465
rect 895 -505 905 -475
rect 935 -505 960 -475
rect 990 -505 1000 -475
rect 895 -515 1000 -505
rect 1145 -475 1250 -465
rect 1145 -505 1155 -475
rect 1185 -505 1210 -475
rect 1240 -505 1250 -475
rect 1145 -515 1250 -505
rect 1395 -475 1500 -465
rect 1395 -505 1405 -475
rect 1435 -505 1460 -475
rect 1490 -505 1500 -475
rect 1395 -515 1500 -505
rect -105 -670 -65 -630
rect -105 -690 -95 -670
rect -75 -690 -65 -670
rect -105 -730 -65 -690
rect -40 -670 0 -515
rect 470 -570 1425 -550
rect 470 -630 490 -570
rect 655 -610 1310 -590
rect 655 -630 675 -610
rect 905 -630 925 -610
rect 1155 -630 1175 -610
rect -40 -690 -30 -670
rect -10 -690 0 -670
rect -40 -730 0 -690
rect 145 -670 185 -630
rect 145 -690 155 -670
rect 175 -690 185 -670
rect 145 -730 185 -690
rect 210 -670 250 -630
rect 395 -670 435 -630
rect 210 -690 220 -670
rect 240 -690 405 -670
rect 425 -690 435 -670
rect 210 -730 250 -690
rect 395 -730 435 -690
rect 460 -670 500 -630
rect 460 -690 470 -670
rect 490 -690 500 -670
rect 460 -730 500 -690
rect 645 -670 685 -630
rect 645 -690 655 -670
rect 675 -690 685 -670
rect 645 -730 685 -690
rect 710 -670 750 -630
rect 710 -690 720 -670
rect 740 -690 750 -670
rect 710 -730 750 -690
rect 895 -670 935 -630
rect 895 -690 905 -670
rect 925 -690 935 -670
rect 895 -730 935 -690
rect 960 -670 1000 -630
rect 960 -690 970 -670
rect 990 -690 1000 -670
rect 960 -730 1000 -690
rect 1145 -670 1185 -630
rect 1145 -690 1155 -670
rect 1175 -690 1185 -670
rect 1145 -730 1185 -690
rect 1210 -670 1250 -630
rect 1210 -690 1220 -670
rect 1240 -690 1250 -670
rect 1210 -730 1250 -690
rect -95 -790 -75 -730
rect 155 -750 175 -730
rect 655 -750 675 -730
rect 155 -770 675 -750
rect 720 -750 740 -730
rect 970 -750 990 -730
rect 1220 -750 1240 -730
rect 720 -770 1240 -750
rect 720 -790 740 -770
rect 1290 -790 1310 -610
rect 1405 -630 1425 -570
rect 1395 -670 1435 -630
rect 1395 -690 1405 -670
rect 1425 -690 1435 -670
rect 1395 -730 1435 -690
rect 1460 -670 1500 -515
rect 1460 -690 1470 -670
rect 1490 -690 1500 -670
rect 1460 -730 1500 -690
rect -95 -810 740 -790
rect 775 -810 1310 -790
rect -170 -835 -125 -820
rect 775 -835 795 -810
rect -170 -855 -155 -835
rect -135 -855 795 -835
rect 905 -855 1425 -835
rect -170 -870 -125 -855
rect -95 -880 -75 -855
rect 155 -880 175 -855
rect 905 -880 925 -855
rect 1155 -880 1175 -855
rect 1405 -880 1425 -855
rect -105 -970 -65 -880
rect -105 -990 -95 -970
rect -75 -990 -65 -970
rect -105 -1080 -65 -990
rect -40 -970 0 -880
rect -40 -990 -30 -970
rect -10 -990 0 -970
rect -40 -1080 0 -990
rect 145 -970 185 -880
rect 145 -990 155 -970
rect 175 -990 185 -970
rect 145 -1080 185 -990
rect 210 -970 250 -880
rect 395 -970 435 -880
rect 210 -990 220 -970
rect 240 -990 405 -970
rect 425 -990 435 -970
rect 210 -1080 250 -990
rect 395 -1080 435 -990
rect 460 -970 500 -880
rect 645 -970 685 -880
rect 460 -990 470 -970
rect 490 -990 655 -970
rect 675 -990 685 -970
rect 460 -1080 500 -990
rect 645 -1080 685 -990
rect 710 -970 750 -880
rect 895 -970 935 -880
rect 710 -990 720 -970
rect 740 -990 905 -970
rect 925 -990 935 -970
rect 710 -1080 750 -990
rect 895 -1080 935 -990
rect 960 -970 1000 -880
rect 960 -990 970 -970
rect 990 -990 1000 -970
rect 960 -1080 1000 -990
rect 1145 -970 1185 -880
rect 1145 -990 1155 -970
rect 1175 -990 1185 -970
rect 1145 -1080 1185 -990
rect 1210 -970 1250 -880
rect 1210 -990 1220 -970
rect 1240 -990 1250 -970
rect 1210 -1080 1250 -990
rect 1395 -970 1435 -880
rect 1395 -990 1405 -970
rect 1425 -990 1435 -970
rect 1395 -1080 1435 -990
rect 1460 -970 1500 -880
rect 1460 -990 1470 -970
rect 1490 -990 1500 -970
rect 1460 -1080 1500 -990
rect -30 -1100 -10 -1080
rect 720 -1100 740 -1080
rect -30 -1120 740 -1100
rect 970 -1100 990 -1080
rect 1220 -1100 1240 -1080
rect 1470 -1100 1490 -1080
rect 970 -1120 1490 -1100
rect 1460 -1140 1490 -1120
rect -105 -1150 0 -1140
rect -105 -1180 -95 -1150
rect -65 -1180 -40 -1150
rect -10 -1180 0 -1150
rect -105 -1190 0 -1180
rect 145 -1150 250 -1140
rect 145 -1180 155 -1150
rect 185 -1180 210 -1150
rect 240 -1180 250 -1150
rect 145 -1190 250 -1180
rect 395 -1150 500 -1140
rect 395 -1180 405 -1150
rect 435 -1180 460 -1150
rect 490 -1180 500 -1150
rect 395 -1190 500 -1180
rect 645 -1150 750 -1140
rect 645 -1180 655 -1150
rect 685 -1180 710 -1150
rect 740 -1180 750 -1150
rect 645 -1190 750 -1180
rect 895 -1150 1000 -1140
rect 895 -1180 905 -1150
rect 935 -1180 960 -1150
rect 990 -1180 1000 -1150
rect 895 -1190 1000 -1180
rect 1145 -1150 1250 -1140
rect 1145 -1180 1155 -1150
rect 1185 -1180 1210 -1150
rect 1240 -1180 1250 -1150
rect 1145 -1190 1250 -1180
rect 1395 -1150 1500 -1140
rect 1395 -1180 1405 -1150
rect 1435 -1180 1460 -1150
rect 1490 -1180 1500 -1150
rect 1395 -1190 1500 -1180
<< viali >>
rect -95 125 -65 155
rect -40 125 -10 155
rect 155 125 185 155
rect 210 125 240 155
rect 405 125 435 155
rect 460 125 490 155
rect 655 125 685 155
rect 710 125 740 155
rect 905 125 935 155
rect 960 125 990 155
rect 1155 125 1185 155
rect 1210 125 1240 155
rect 1405 125 1435 155
rect 1460 125 1490 155
rect 265 -255 285 -235
rect 1140 -200 1160 -180
rect 1390 -200 1410 -180
rect 1475 -185 1495 -165
rect 1225 -265 1245 -245
rect -95 -505 -65 -475
rect -40 -505 -10 -475
rect 155 -505 185 -475
rect 210 -505 240 -475
rect 405 -505 435 -475
rect 460 -505 490 -475
rect 655 -505 685 -475
rect 710 -505 740 -475
rect 905 -505 935 -475
rect 960 -505 990 -475
rect 1155 -505 1185 -475
rect 1210 -505 1240 -475
rect 1405 -505 1435 -475
rect 1460 -505 1490 -475
rect -155 -855 -135 -835
rect -95 -1180 -65 -1150
rect -40 -1180 -10 -1150
rect 155 -1180 185 -1150
rect 210 -1180 240 -1150
rect 405 -1180 435 -1150
rect 460 -1180 490 -1150
rect 655 -1180 685 -1150
rect 710 -1180 740 -1150
rect 905 -1180 935 -1150
rect 960 -1180 990 -1150
rect 1155 -1180 1185 -1150
rect 1210 -1180 1240 -1150
rect 1405 -1180 1435 -1150
rect 1460 -1180 1490 -1150
<< metal1 >>
rect -250 155 1660 165
rect -250 125 -95 155
rect -65 125 -40 155
rect -10 125 155 155
rect 185 125 210 155
rect 240 125 405 155
rect 435 125 460 155
rect 490 125 655 155
rect 685 125 710 155
rect 740 125 905 155
rect 935 125 960 155
rect 990 125 1155 155
rect 1185 125 1210 155
rect 1240 125 1405 155
rect 1435 125 1460 155
rect 1490 125 1660 155
rect -250 115 1660 125
rect 1500 -155 1660 -150
rect 1465 -165 1660 -155
rect 1040 -180 1180 -170
rect -245 -235 295 -185
rect 1040 -200 1140 -180
rect 1160 -200 1180 -180
rect 1040 -210 1180 -200
rect 1290 -180 1430 -170
rect 1290 -200 1390 -180
rect 1410 -200 1430 -180
rect 1465 -185 1475 -165
rect 1495 -185 1660 -165
rect 1465 -200 1660 -185
rect 1290 -210 1430 -200
rect 1250 -230 1660 -225
rect 255 -255 265 -235
rect 285 -255 295 -235
rect 255 -265 295 -255
rect 1215 -245 1660 -230
rect 1215 -265 1225 -245
rect 1245 -265 1660 -245
rect 1215 -275 1660 -265
rect -250 -475 1660 -465
rect -250 -505 -95 -475
rect -65 -505 -40 -475
rect -10 -505 155 -475
rect 185 -505 210 -475
rect 240 -505 405 -475
rect 435 -505 460 -475
rect 490 -505 655 -475
rect 685 -505 710 -475
rect 740 -505 905 -475
rect 935 -505 960 -475
rect 990 -505 1155 -475
rect 1185 -505 1210 -475
rect 1240 -505 1405 -475
rect 1435 -505 1460 -475
rect 1490 -505 1660 -475
rect -250 -515 1660 -505
rect -250 -835 -110 -820
rect -250 -855 -155 -835
rect -135 -855 -110 -835
rect -250 -870 -110 -855
rect -250 -1150 1660 -1140
rect -250 -1180 -95 -1150
rect -65 -1180 -40 -1150
rect -10 -1180 155 -1150
rect 185 -1180 210 -1150
rect 240 -1180 405 -1150
rect 435 -1180 460 -1150
rect 490 -1180 655 -1150
rect 685 -1180 710 -1150
rect 740 -1180 905 -1150
rect 935 -1180 960 -1150
rect 990 -1180 1155 -1150
rect 1185 -1180 1210 -1150
rect 1240 -1180 1405 -1150
rect 1435 -1180 1460 -1150
rect 1490 -1180 1660 -1150
rect -250 -1190 1660 -1180
<< labels >>
rlabel metal1 -250 115 -250 165 3 vdd
rlabel metal1 -250 -1190 -250 -1140 3 gnd
rlabel metal1 -250 -1190 -250 -1140 3 vdd
rlabel metal1 -250 -515 -250 -465 3 gnd
rlabel metal1 -245 -235 -245 -185 1 cout_comp
rlabel metal1 1040 -210 1040 -170 1 cout_comp
rlabel metal1 1290 -210 1290 -170 1 sum_comp
rlabel metal1 1660 -200 1660 -150 7 sum
rlabel metal1 1660 -275 1660 -225 7 cout
rlabel metal1 -250 -870 -250 -820 3 sum_comp
rlabel poly -60 65 -45 65 1 b
rlabel poly 190 65 205 65 1 a
rlabel poly 440 65 455 65 1 a
rlabel poly 690 65 705 65 1 b
rlabel poly 940 65 955 65 1 cin
rlabel poly -60 -1095 -45 -1095 1 cout_comp
rlabel poly 190 -1095 205 -1095 1 a
rlabel poly 440 -1095 455 -1095 1 b
rlabel poly 690 -1095 705 -1095 1 cin
rlabel poly 940 -1095 955 -1095 1 b
rlabel poly 1190 -1095 1205 -1095 1 a
rlabel poly 1440 -1095 1455 -1095 1 cin
<< end >>
